//package where all the classes are included

`include "seq_item.sv"
`include "reg_pkg.sv"
`include "reg_apb_adapter.sv"
`include "base_seq.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "environment.sv"

